`timescale 1ns/1ps

module dff (
    input  logic clk,
    input  logic rst,
    input  logic d,
    output logic q
);

always_ff @(posedge clk) begin
    if (rst)
        q <= 1'b0;
    else
        q <= d;
end

endmodule
